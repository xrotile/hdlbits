module top_module (
    input in,
    output out);
	assign out = in;
endmodule

